`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/23/2025 02:49:58 PM
// Design Name: 
// Module Name: warning_system_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module warning_system_tb(

    );
    
 

	//regs for inputs
	//SB, DOOR, KEY, BRK, PARK, HOOD, BAT_OK, AIB_OK, TMP_OK, PASS_OCC, SB_P, TRUNK, PBRK, SRV
	reg [0:13] i;
	//wires for outputs
	wire START_PERMIT, CHIME, WARN_PRI2, WARN_PRI1, SEAT_WARN, DOOR_WARN, HOOD_WARN, TRUNK_WARN, BAT_WARN, AIRBAG_WARN, TEMP_WARN;
	
	//instantiate module to test
	warning_system uut(.i({i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], i[4], i[3], i[2], i[1], i[0]}),
					.o({WARN_PRI1, TEMP_WARN, AIRBAG_WARN, BAT_WARN, TRUNK_WARN, HOOD_WARN, DOOR_WARN, SEAT_WARN, CHIME, START_PERMIT, WARN_PRI2}));
	//WARN_PRI1, TEMP_WARN, AIRBAG_WARN, BAT_WARN, TRUNK_WARN, HOOD_WARN, DOOR_WARN, SEAT_WARN, CHIME, START_PERMIT, WARN_PRI2
	//test cases
	initial begin
		i = 14'b0;
		//car can start normally
		i[2]=1; i[3]=1; i[4]=1; i[6]=1; i[7]=1; i[8]=1;
		#10;
		
		//car cannot start because no key
		i[2] = 0;
		#10;
		
		i = 14'b0;
		//car can start to be serviced
		i[2]=1; i[3]=1; i[4]=1; i[6]=0; i[7]=0; i[8]=0; i[13]=1;
		#10;
		
		i = 14'b0;
		//driver seatbelt unbuckled
		i[0] = 0;
		#10;
		
		i = 14'b0;
		//passenger is present and seatbelt unbuckled
		i[9] = 1; i[10] = 0;
		#10;
		
		i = 14'b0;
		//door is open
		i[1]=0;
		#10;
		
		i = 14'b0;
		//hood is open
		i[5]=0;
		#10;
		
		i = 14'b0;
		//trunk is open
		i[11]=0;
		#10;
		
		i = 14'b0;
		//battery not okay
		i[6]=0;
		#10;
		
		i = 14'b0;
		//airbag not okay
		i[7]=0;
		#10;
		
		i = 14'b0;
		//coolant temp not okay
		i[8]=0;
		#10;
		
		i = 14'b0;
		//parking brake on
		i[12]=1;
		#10;
		$stop;




	end
endmodule
   
